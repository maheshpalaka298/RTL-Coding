`timescale 1ns / 1ps

//Author Name : Mahesh Palaka
//Project Name: Parallel-in-Parallel-out shift Register

module pipo_reg(clk,clear,d,q);

  input clk,clear;

  output reg [3:0]  q;
  input [3:0] d;


  always @(posedge clk )
    begin
      if (clear)
        q <= 4'b0000;
      else
        q <= d;
    end
endmodule`timescale 1ns / 1ps

//Author Name : Mahesh Palaka
//Project Name: Bi-Driectional shift Register

module bidirectional_reg  #(parameter MSB=4) (input d,                      // Declare input for data to the first flop in the shift register
                                        input clk,                    // Declare input for clock to all flops in the shift register
                                        input en,                     // Declare input for enable to switch the shift register on/off
                                        input dir,                    // Declare input to shift in either left or right direction
                                        input rstn,                   // Declare input to reset the register to a default value
                                        output reg [MSB-1:0] out);    // Declare output to read out the current value of all flops in this register


   always @ (posedge clk)
      if (!rstn)
         out <= 0;
      else begin
         if (en)
            case (dir)
               0 :  out <= {out[MSB-2:0], d};
               1 :  out <= {d, out[MSB-1:1]};
            endcase
         else
            out <= out;
      end
endmodule
